module cons(output wire [31:0] cero, cuatro, menos_cuatro);
	assign cero = 32'sd0;
	assign cuatro = 32'sd4;
	assign menos_cuatro = -32'sd4;
endmodule